LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.ALL;

ENTITY GammaCorrection IS
  PORT (
    input   : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    output  : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END ENTITY;

ARCHITECTURE arch OF GammaCorrection IS
  BEGIN
  PROCESS (input) IS
    BEGIN
      CASE input IS      
        WHEN "00000000" => output <= "00000000";
        WHEN "00000001" => output <= "00000000";
        WHEN "00000010" => output <= "00000000";
        WHEN "00000011" => output <= "00000000";
        WHEN "00000100" => output <= "00000000";
        WHEN "00000101" => output <= "00000000";
        WHEN "00000110" => output <= "00000000";
        WHEN "00000111" => output <= "00000000";
        WHEN "00001000" => output <= "00000000";
        WHEN "00001001" => output <= "00000000";
        WHEN "00001010" => output <= "00000000";
        WHEN "00001011" => output <= "00000000";
        WHEN "00001100" => output <= "00000000";
        WHEN "00001101" => output <= "00000000";
        WHEN "00001110" => output <= "00000000";
        WHEN "00001111" => output <= "00000000";
        WHEN "00010000" => output <= "00000000";
        WHEN "00010001" => output <= "00000000";
        WHEN "00010010" => output <= "00000000";
        WHEN "00010011" => output <= "00000000";
        WHEN "00010100" => output <= "00000000";
        WHEN "00010101" => output <= "00000000";
        WHEN "00010110" => output <= "00000000";
        WHEN "00010111" => output <= "00000000";
        WHEN "00011000" => output <= "00000000";
        WHEN "00011001" => output <= "00000000";
        WHEN "00011010" => output <= "00000000";
        WHEN "00011011" => output <= "00000000";
        WHEN "00011100" => output <= "00000000";
        WHEN "00011101" => output <= "00000000";
        WHEN "00011110" => output <= "00000000";
        WHEN "00011111" => output <= "00000000";
        WHEN "00100000" => output <= "00000000";
        WHEN "00100001" => output <= "00000000";
        WHEN "00100010" => output <= "00000000";
        WHEN "00100011" => output <= "00000000";
        WHEN "00100100" => output <= "00000000";
        WHEN "00100101" => output <= "00000000";
        WHEN "00100110" => output <= "00000000";
        WHEN "00100111" => output <= "00000000";
        WHEN "00101000" => output <= "00000000";
        WHEN "00101001" => output <= "00000000";
        WHEN "00101010" => output <= "00000000";
        WHEN "00101011" => output <= "00000000";
        WHEN "00101100" => output <= "00000000";
        WHEN "00101101" => output <= "00000000";
        WHEN "00101110" => output <= "00000000";
        WHEN "00101111" => output <= "00000000";
        WHEN "00110000" => output <= "00000000";
        WHEN "00110001" => output <= "00000001";
        WHEN "00110010" => output <= "00000001";
        WHEN "00110011" => output <= "00000001";
        WHEN "00110100" => output <= "00000001";
        WHEN "00110101" => output <= "00000001";
        WHEN "00110110" => output <= "00000001";
        WHEN "00110111" => output <= "00000001";
        WHEN "00111000" => output <= "00000001";
        WHEN "00111001" => output <= "00000001";
        WHEN "00111010" => output <= "00000001";
        WHEN "00111011" => output <= "00000001";
        WHEN "00111100" => output <= "00000010";
        WHEN "00111101" => output <= "00000010";
        WHEN "00111110" => output <= "00000010";
        WHEN "00111111" => output <= "00000010";
        WHEN "01000000" => output <= "00000010";
        WHEN "01000001" => output <= "00000010";
        WHEN "01000010" => output <= "00000010";
        WHEN "01000011" => output <= "00000010";
        WHEN "01000100" => output <= "00000011";
        WHEN "01000101" => output <= "00000011";
        WHEN "01000110" => output <= "00000011";
        WHEN "01000111" => output <= "00000011";
        WHEN "01001000" => output <= "00000011";
        WHEN "01001001" => output <= "00000011";
        WHEN "01001010" => output <= "00000100";
        WHEN "01001011" => output <= "00000100";
        WHEN "01001100" => output <= "00000100";
        WHEN "01001101" => output <= "00000100";
        WHEN "01001110" => output <= "00000100";
        WHEN "01001111" => output <= "00000101";
        WHEN "01010000" => output <= "00000101";
        WHEN "01010001" => output <= "00000101";
        WHEN "01010010" => output <= "00000101";
        WHEN "01010011" => output <= "00000110";
        WHEN "01010100" => output <= "00000110";
        WHEN "01010101" => output <= "00000110";
        WHEN "01010110" => output <= "00000110";
        WHEN "01010111" => output <= "00000111";
        WHEN "01011000" => output <= "00000111";
        WHEN "01011001" => output <= "00000111";
        WHEN "01011010" => output <= "00000111";
        WHEN "01011011" => output <= "00001000";
        WHEN "01011100" => output <= "00001000";
        WHEN "01011101" => output <= "00001000";
        WHEN "01011110" => output <= "00001001";
        WHEN "01011111" => output <= "00001001";
        WHEN "01100000" => output <= "00001001";
        WHEN "01100001" => output <= "00001010";
        WHEN "01100010" => output <= "00001010";
        WHEN "01100011" => output <= "00001010";
        WHEN "01100100" => output <= "00001011";
        WHEN "01100101" => output <= "00001011";
        WHEN "01100110" => output <= "00001100";
        WHEN "01100111" => output <= "00001100";
        WHEN "01101000" => output <= "00001100";
        WHEN "01101001" => output <= "00001101";
        WHEN "01101010" => output <= "00001101";
        WHEN "01101011" => output <= "00001110";
        WHEN "01101100" => output <= "00001110";
        WHEN "01101101" => output <= "00001111";
        WHEN "01101110" => output <= "00001111";
        WHEN "01101111" => output <= "00001111";
        WHEN "01110000" => output <= "00010000";
        WHEN "01110001" => output <= "00010000";
        WHEN "01110010" => output <= "00010001";
        WHEN "01110011" => output <= "00010001";
        WHEN "01110100" => output <= "00010010";
        WHEN "01110101" => output <= "00010010";
        WHEN "01110110" => output <= "00010011";
        WHEN "01110111" => output <= "00010100";
        WHEN "01111000" => output <= "00010100";
        WHEN "01111001" => output <= "00010101";
        WHEN "01111010" => output <= "00010101";
        WHEN "01111011" => output <= "00010110";
        WHEN "01111100" => output <= "00010111";
        WHEN "01111101" => output <= "00010111";
        WHEN "01111110" => output <= "00011000";
        WHEN "01111111" => output <= "00011000";
        WHEN "10000000" => output <= "00011001";
        WHEN "10000001" => output <= "00011010";
        WHEN "10000010" => output <= "00011010";
        WHEN "10000011" => output <= "00011011";
        WHEN "10000100" => output <= "00011100";
        WHEN "10000101" => output <= "00011101";
        WHEN "10000110" => output <= "00011101";
        WHEN "10000111" => output <= "00011110";
        WHEN "10001000" => output <= "00011111";
        WHEN "10001001" => output <= "00100000";
        WHEN "10001010" => output <= "00100000";
        WHEN "10001011" => output <= "00100001";
        WHEN "10001100" => output <= "00100010";
        WHEN "10001101" => output <= "00100011";
        WHEN "10001110" => output <= "00100100";
        WHEN "10001111" => output <= "00100101";
        WHEN "10010000" => output <= "00100101";
        WHEN "10010001" => output <= "00100110";
        WHEN "10010010" => output <= "00100111";
        WHEN "10010011" => output <= "00101000";
        WHEN "10010100" => output <= "00101001";
        WHEN "10010101" => output <= "00101010";
        WHEN "10010110" => output <= "00101011";
        WHEN "10010111" => output <= "00101100";
        WHEN "10011000" => output <= "00101101";
        WHEN "10011001" => output <= "00101110";
        WHEN "10011010" => output <= "00101111";
        WHEN "10011011" => output <= "00110000";
        WHEN "10011100" => output <= "00110001";
        WHEN "10011101" => output <= "00110010";
        WHEN "10011110" => output <= "00110011";
        WHEN "10011111" => output <= "00110100";
        WHEN "10100000" => output <= "00110101";
        WHEN "10100001" => output <= "00110111";
        WHEN "10100010" => output <= "00111000";
        WHEN "10100011" => output <= "00111001";
        WHEN "10100100" => output <= "00111010";
        WHEN "10100101" => output <= "00111011";
        WHEN "10100110" => output <= "00111100";
        WHEN "10100111" => output <= "00111110";
        WHEN "10101000" => output <= "00111111";
        WHEN "10101001" => output <= "01000000";
        WHEN "10101010" => output <= "01000010";
        WHEN "10101011" => output <= "01000011";
        WHEN "10101100" => output <= "01000100";
        WHEN "10101101" => output <= "01000101";
        WHEN "10101110" => output <= "01000111";
        WHEN "10101111" => output <= "01001000";
        WHEN "10110000" => output <= "01001010";
        WHEN "10110001" => output <= "01001011";
        WHEN "10110010" => output <= "01001100";
        WHEN "10110011" => output <= "01001110";
        WHEN "10110100" => output <= "01001111";
        WHEN "10110101" => output <= "01010001";
        WHEN "10110110" => output <= "01010010";
        WHEN "10110111" => output <= "01010100";
        WHEN "10111000" => output <= "01010101";
        WHEN "10111001" => output <= "01010111";
        WHEN "10111010" => output <= "01011001";
        WHEN "10111011" => output <= "01011010";
        WHEN "10111100" => output <= "01011100";
        WHEN "10111101" => output <= "01011101";
        WHEN "10111110" => output <= "01011111";
        WHEN "10111111" => output <= "01100001";
        WHEN "11000000" => output <= "01100011";
        WHEN "11000001" => output <= "01100100";
        WHEN "11000010" => output <= "01100110";
        WHEN "11000011" => output <= "01101000";
        WHEN "11000100" => output <= "01101010";
        WHEN "11000101" => output <= "01101011";
        WHEN "11000110" => output <= "01101101";
        WHEN "11000111" => output <= "01101111";
        WHEN "11001000" => output <= "01110001";
        WHEN "11001001" => output <= "01110011";
        WHEN "11001010" => output <= "01110101";
        WHEN "11001011" => output <= "01110111";
        WHEN "11001100" => output <= "01111001";
        WHEN "11001101" => output <= "01111011";
        WHEN "11001110" => output <= "01111101";
        WHEN "11001111" => output <= "01111111";
        WHEN "11010000" => output <= "10000001";
        WHEN "11010001" => output <= "10000011";
        WHEN "11010010" => output <= "10000101";
        WHEN "11010011" => output <= "10000111";
        WHEN "11010100" => output <= "10001001";
        WHEN "11010101" => output <= "10001011";
        WHEN "11010110" => output <= "10001110";
        WHEN "11010111" => output <= "10010000";
        WHEN "11011000" => output <= "10010010";
        WHEN "11011001" => output <= "10010100";
        WHEN "11011010" => output <= "10010111";
        WHEN "11011011" => output <= "10011001";
        WHEN "11011100" => output <= "10011011";
        WHEN "11011101" => output <= "10011110";
        WHEN "11011110" => output <= "10100000";
        WHEN "11011111" => output <= "10100011";
        WHEN "11100000" => output <= "10100101";
        WHEN "11100001" => output <= "10101000";
        WHEN "11100010" => output <= "10101010";
        WHEN "11100011" => output <= "10101101";
        WHEN "11100100" => output <= "10101111";
        WHEN "11100101" => output <= "10110010";
        WHEN "11100110" => output <= "10110100";
        WHEN "11100111" => output <= "10110111";
        WHEN "11101000" => output <= "10111010";
        WHEN "11101001" => output <= "10111100";
        WHEN "11101010" => output <= "10111111";
        WHEN "11101011" => output <= "11000010";
        WHEN "11101100" => output <= "11000100";
        WHEN "11101101" => output <= "11000111";
        WHEN "11101110" => output <= "11001010";
        WHEN "11101111" => output <= "11001101";
        WHEN "11110000" => output <= "11010000";
        WHEN "11110001" => output <= "11010011";
        WHEN "11110010" => output <= "11010110";
        WHEN "11110011" => output <= "11011001";
        WHEN "11110100" => output <= "11011100";
        WHEN "11110101" => output <= "11011111";
        WHEN "11110110" => output <= "11100010";
        WHEN "11110111" => output <= "11100101";
        WHEN "11111000" => output <= "11101000";
        WHEN "11111001" => output <= "11101011";
        WHEN "11111010" => output <= "11101110";
        WHEN "11111011" => output <= "11110001";
        WHEN "11111100" => output <= "11110101";
        WHEN "11111101" => output <= "11111000";
        WHEN "11111110" => output <= "11111011";
        WHEN "11111111" => output <= "11111111";
        WHEN OTHERS => output <= input;
      END CASE;
  END PROCESS;
END ARCHITECTURE; 